//This is tb_memory, get input from FPGA, and store here

`timescale 1ns / 1ps

module tb_memory;

endmodule
