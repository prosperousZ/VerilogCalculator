//This is tb_datapath file


`timescale 1ns / 1ps

module tb_datapath;



endmodule
