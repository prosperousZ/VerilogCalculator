//This is tb_io_interface file

`timescale 1ns / 1ps

module tb_io_interface;

endmodule
