//This is io_vga file, display on screen, i am not sure if we want to diplay
//on the LCD screen, or just display on FPGA, may not need this file


module io_vga();


endmodule
