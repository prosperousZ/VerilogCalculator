
//////////////////////////////////////////////////////////////////////////////////
// Module Name:		io_interface
// Description: 	Module to interface between the chip and the FPGA
//
// Dependencies: 	
//
// Comments: 		
//
//////////////////////////////////////////////////////////////////////////////////
module io_interface();

endmodule
