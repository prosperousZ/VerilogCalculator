//this is test bench of finalProject
`timescale 1ns / 1ps


module tb_finalProject;

endmodule
