//////////////////////////////////////////////////////////////////////////////////
// Module Name:		regfile
// Description: 	
//
// Dependencies: 	
//
// Comments: 		
//
//////////////////////////////////////////////////////////////////////////////////
module regfile();

endmodule
