// This is the regfile


module regfile();

endmodule
