
//This is io_interface file， interface between chip and FPGA

module io_interface();

endmodule
