//This is tb_alu file
`timescale 1ns / 1ps

module tb_alu;

endmodule
