//This memory file, to store previous output

module memory();


endmodule
