//This is tb_processor file

`timescale 1ns / 1ps

module tb_processor;

endmodule
